class driver;

endclass

