module dut_top (
    input   clk
);
    initial begin
        $display("dut_top module");
    end
endmodule
